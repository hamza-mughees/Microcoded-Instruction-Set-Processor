library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity control_memory is
	port (
		in_car : in std_logic_vector (7 downto 0);
		mw, mm, rw, md : out std_logic;
		fs : out std_logic_vector (4 downto 0);
		mb, tb, ta, td, pl, pi, il, mc : out std_logic;
		ms : out std_logic_vector (2 downto 0);
		na : out std_logic_vector (7 downto 0)
	);
end control_memory;

architecture dataflow of control_memory is
	type mem_array is array (0 to 255) of std_logic_vector (27 downto 0);
begin
	memory_m: process (in_car)
		variable control_mem : mem_array := (
			-- 0
			x"fffffff",	-- 0
			x"0000000",	-- 1
			x"aaaaaaa",	-- 2
			x"0000000",	-- 3
			x"bbbbbbb",	-- 4
			x"0000000",	-- 5
			x"ccccccc",	-- 6
			x"0000000",	-- 7
			x"ddddddd",	-- 8
			x"0000000",	-- 9
			x"1111111",	-- a
			x"0000000",	-- b
			x"2222222",	-- c
			x"0000000",	-- d
			x"3333333",	-- e
			x"0000000",	-- f
			
			-- 1
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- 2
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- 3
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- 4
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- 5
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- 6
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- 7
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- 8
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- 9
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- a
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- b
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- c
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- d 
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- e 
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
			
			-- f
			x"0000000",	-- 0
			x"0000000",	-- 1
			x"0000000",	-- 2
			x"0000000",	-- 3
			x"0000000",	-- 4
			x"0000000",	-- 5
			x"0000000",	-- 6
			x"0000000",	-- 7
			x"0000000",	-- 8
			x"0000000",	-- 9
			x"0000000",	-- a
			x"0000000",	-- b
			x"0000000",	-- c
			x"0000000",	-- d
			x"0000000",	-- e
			x"0000000",	-- f
		);
	
		variable addr : integer;
		variable control_out : std_logic_vector (27 downto 0);
	begin
		addr := conv_integer(in_car);
		control_out := control_mem(addr);
		mw <= control_out(0);
		mm <= control_out(1);
		rw <= control_out(2);
		md <= control_out(3);
		fs <= control_out(8 downto 4);
		mb <= control_out(9);
		tb <= control_out(10);
		ta <= control_out(11);
		td <= control_out(12);
		pl <= control_out(13);
		pi <= control_out(14);
		il <= control_out(15);
		mc <= control_out(16);
		ns <= control_out(19 downto 17);
		na <= control_out(27 downto 20);
	end process;
end dataflow;