library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity external_memory is
	port (
		address, data_to_write : in std_logic_vector (15 downto 0);
		write_to_mem, Clk : in std_logic;
		data_to_read : out std_logic_vector (15 downto 0)
	);
end external_memory;

architecture dataflow of external_memory is
	type mem_array is array (0 to 511) of std_logic_vector (15 downto 0);
begin
	memory: process (address, data_to_write, Clk)
		variable data_mem : mem_array := (
			x"0abc", x"0123", x"05ad", x"0fd3",
			x"0110", x"0efe", x"0f75", x"05b6",
			x"0c4a", x"09ab", x"0cf9", x"088a",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
			x"0000", x"0000", x"0000", x"0000",
		);
		
		variable addr : integer;
	begin
		addr := conv_integer(unsigned(address(8 downto 0)));
		-- ^ least significant 9 bits used to index into array
		if write_to_mem="1" then
			data_mem(addr) := data_to_write;
		else
			data_to_read <= data_mem(addr) after 5ns;
	end process;
end dataflow;